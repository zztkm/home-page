module main

fn hello() string {
	return "Hello!"
}

fn main() {
	println(hello())
}
